// system_acl_iface.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module system_acl_iface (
		output wire [1:0]   acl_internal_memorg_kernel_mode,         //       acl_internal_memorg_kernel.mode
		output wire         acl_kernel_clk_kernel_pll_locked_export, // acl_kernel_clk_kernel_pll_locked.export
		input  wire         config_clk_clk,                          //                       config_clk.clk
		input  wire         reset_n,                                 //                     global_reset.reset_n
		output wire         kernel_clk_clk,                          //                       kernel_clk.clk
		output wire         kernel_clk2x_clk,                        //                     kernel_clk2x.clk
		output wire         kernel_clk_snoop_clk,                    //                 kernel_clk_snoop.clk
		input  wire         kernel_cra_waitrequest,                  //                       kernel_cra.waitrequest
		input  wire [63:0]  kernel_cra_readdata,                     //                                 .readdata
		input  wire         kernel_cra_readdatavalid,                //                                 .readdatavalid
		output wire [0:0]   kernel_cra_burstcount,                   //                                 .burstcount
		output wire [63:0]  kernel_cra_writedata,                    //                                 .writedata
		output wire [29:0]  kernel_cra_address,                      //                                 .address
		output wire         kernel_cra_write,                        //                                 .write
		output wire         kernel_cra_read,                         //                                 .read
		output wire [7:0]   kernel_cra_byteenable,                   //                                 .byteenable
		output wire         kernel_cra_debugaccess,                  //                                 .debugaccess
		input  wire [0:0]   kernel_irq_irq,                          //                       kernel_irq.irq
		output wire         kernel_mem0_waitrequest,                 //                      kernel_mem0.waitrequest
		output wire [255:0] kernel_mem0_readdata,                    //                                 .readdata
		output wire         kernel_mem0_readdatavalid,               //                                 .readdatavalid
		input  wire [4:0]   kernel_mem0_burstcount,                  //                                 .burstcount
		input  wire [255:0] kernel_mem0_writedata,                   //                                 .writedata
		input  wire [24:0]  kernel_mem0_address,                     //                                 .address
		input  wire         kernel_mem0_write,                       //                                 .write
		input  wire         kernel_mem0_read,                        //                                 .read
		input  wire [31:0]  kernel_mem0_byteenable,                  //                                 .byteenable
		input  wire         kernel_mem0_debugaccess,                 //                                 .debugaccess
		input  wire         kernel_pll_refclk_clk,                   //                kernel_pll_refclk.clk
		output wire         kernel_reset_reset_n,                    //                     kernel_reset.reset_n
		output wire [14:0]  memory_mem_a,                            //                           memory.mem_a
		output wire [2:0]   memory_mem_ba,                           //                                 .mem_ba
		output wire         memory_mem_ck,                           //                                 .mem_ck
		output wire         memory_mem_ck_n,                         //                                 .mem_ck_n
		output wire         memory_mem_cke,                          //                                 .mem_cke
		output wire         memory_mem_cs_n,                         //                                 .mem_cs_n
		output wire         memory_mem_ras_n,                        //                                 .mem_ras_n
		output wire         memory_mem_cas_n,                        //                                 .mem_cas_n
		output wire         memory_mem_we_n,                         //                                 .mem_we_n
		output wire         memory_mem_reset_n,                      //                                 .mem_reset_n
		inout  wire [31:0]  memory_mem_dq,                           //                                 .mem_dq
		inout  wire [3:0]   memory_mem_dqs,                          //                                 .mem_dqs
		inout  wire [3:0]   memory_mem_dqs_n,                        //                                 .mem_dqs_n
		output wire         memory_mem_odt,                          //                                 .mem_odt
		output wire [3:0]   memory_mem_dm,                           //                                 .mem_dm
		input  wire         memory_oct_rzqin,                        //                                 .oct_rzqin
		output wire         peripheral_hps_io_emac1_inst_TX_CLK,     //                       peripheral.hps_io_emac1_inst_TX_CLK
		output wire         peripheral_hps_io_emac1_inst_TXD0,       //                                 .hps_io_emac1_inst_TXD0
		output wire         peripheral_hps_io_emac1_inst_TXD1,       //                                 .hps_io_emac1_inst_TXD1
		output wire         peripheral_hps_io_emac1_inst_TXD2,       //                                 .hps_io_emac1_inst_TXD2
		output wire         peripheral_hps_io_emac1_inst_TXD3,       //                                 .hps_io_emac1_inst_TXD3
		input  wire         peripheral_hps_io_emac1_inst_RXD0,       //                                 .hps_io_emac1_inst_RXD0
		inout  wire         peripheral_hps_io_emac1_inst_MDIO,       //                                 .hps_io_emac1_inst_MDIO
		output wire         peripheral_hps_io_emac1_inst_MDC,        //                                 .hps_io_emac1_inst_MDC
		input  wire         peripheral_hps_io_emac1_inst_RX_CTL,     //                                 .hps_io_emac1_inst_RX_CTL
		output wire         peripheral_hps_io_emac1_inst_TX_CTL,     //                                 .hps_io_emac1_inst_TX_CTL
		input  wire         peripheral_hps_io_emac1_inst_RX_CLK,     //                                 .hps_io_emac1_inst_RX_CLK
		input  wire         peripheral_hps_io_emac1_inst_RXD1,       //                                 .hps_io_emac1_inst_RXD1
		input  wire         peripheral_hps_io_emac1_inst_RXD2,       //                                 .hps_io_emac1_inst_RXD2
		input  wire         peripheral_hps_io_emac1_inst_RXD3,       //                                 .hps_io_emac1_inst_RXD3
		inout  wire         peripheral_hps_io_sdio_inst_CMD,         //                                 .hps_io_sdio_inst_CMD
		inout  wire         peripheral_hps_io_sdio_inst_D0,          //                                 .hps_io_sdio_inst_D0
		inout  wire         peripheral_hps_io_sdio_inst_D1,          //                                 .hps_io_sdio_inst_D1
		output wire         peripheral_hps_io_sdio_inst_CLK,         //                                 .hps_io_sdio_inst_CLK
		inout  wire         peripheral_hps_io_sdio_inst_D2,          //                                 .hps_io_sdio_inst_D2
		inout  wire         peripheral_hps_io_sdio_inst_D3,          //                                 .hps_io_sdio_inst_D3
		inout  wire         peripheral_hps_io_usb1_inst_D0,          //                                 .hps_io_usb1_inst_D0
		inout  wire         peripheral_hps_io_usb1_inst_D1,          //                                 .hps_io_usb1_inst_D1
		inout  wire         peripheral_hps_io_usb1_inst_D2,          //                                 .hps_io_usb1_inst_D2
		inout  wire         peripheral_hps_io_usb1_inst_D3,          //                                 .hps_io_usb1_inst_D3
		inout  wire         peripheral_hps_io_usb1_inst_D4,          //                                 .hps_io_usb1_inst_D4
		inout  wire         peripheral_hps_io_usb1_inst_D5,          //                                 .hps_io_usb1_inst_D5
		inout  wire         peripheral_hps_io_usb1_inst_D6,          //                                 .hps_io_usb1_inst_D6
		inout  wire         peripheral_hps_io_usb1_inst_D7,          //                                 .hps_io_usb1_inst_D7
		input  wire         peripheral_hps_io_usb1_inst_CLK,         //                                 .hps_io_usb1_inst_CLK
		output wire         peripheral_hps_io_usb1_inst_STP,         //                                 .hps_io_usb1_inst_STP
		input  wire         peripheral_hps_io_usb1_inst_DIR,         //                                 .hps_io_usb1_inst_DIR
		input  wire         peripheral_hps_io_usb1_inst_NXT,         //                                 .hps_io_usb1_inst_NXT
		input  wire         peripheral_hps_io_uart0_inst_RX,         //                                 .hps_io_uart0_inst_RX
		output wire         peripheral_hps_io_uart0_inst_TX,         //                                 .hps_io_uart0_inst_TX
		inout  wire         peripheral_hps_io_i2c1_inst_SDA,         //                                 .hps_io_i2c1_inst_SDA
		inout  wire         peripheral_hps_io_i2c1_inst_SCL,         //                                 .hps_io_i2c1_inst_SCL
		inout  wire         peripheral_hps_io_gpio_inst_GPIO53       //                                 .hps_io_gpio_inst_GPIO53
	);

	wire          pll_outclk0_clk;                                                             // pll:outclk_0 -> [address_span_extender_kernel:clk, clock_cross_kernel_mem1:m0_clk, hps:f2h_sdram0_clk, mm_interconnect_0:pll_outclk0_clk, mm_interconnect_3:pll_outclk0_clk, rst_controller_001:clk, rst_controller_002:clk]
	wire          address_span_extender_kernel_expanded_master_waitrequest;                    // mm_interconnect_0:address_span_extender_kernel_expanded_master_waitrequest -> address_span_extender_kernel:avm_m0_waitrequest
	wire  [255:0] address_span_extender_kernel_expanded_master_readdata;                       // mm_interconnect_0:address_span_extender_kernel_expanded_master_readdata -> address_span_extender_kernel:avm_m0_readdata
	wire   [31:0] address_span_extender_kernel_expanded_master_address;                        // address_span_extender_kernel:avm_m0_address -> mm_interconnect_0:address_span_extender_kernel_expanded_master_address
	wire          address_span_extender_kernel_expanded_master_read;                           // address_span_extender_kernel:avm_m0_read -> mm_interconnect_0:address_span_extender_kernel_expanded_master_read
	wire   [31:0] address_span_extender_kernel_expanded_master_byteenable;                     // address_span_extender_kernel:avm_m0_byteenable -> mm_interconnect_0:address_span_extender_kernel_expanded_master_byteenable
	wire          address_span_extender_kernel_expanded_master_readdatavalid;                  // mm_interconnect_0:address_span_extender_kernel_expanded_master_readdatavalid -> address_span_extender_kernel:avm_m0_readdatavalid
	wire          address_span_extender_kernel_expanded_master_write;                          // address_span_extender_kernel:avm_m0_write -> mm_interconnect_0:address_span_extender_kernel_expanded_master_write
	wire  [255:0] address_span_extender_kernel_expanded_master_writedata;                      // address_span_extender_kernel:avm_m0_writedata -> mm_interconnect_0:address_span_extender_kernel_expanded_master_writedata
	wire    [4:0] address_span_extender_kernel_expanded_master_burstcount;                     // address_span_extender_kernel:avm_m0_burstcount -> mm_interconnect_0:address_span_extender_kernel_expanded_master_burstcount
	wire  [255:0] mm_interconnect_0_hps_f2h_sdram0_data_readdata;                              // hps:f2h_sdram0_READDATA -> mm_interconnect_0:hps_f2h_sdram0_data_readdata
	wire          mm_interconnect_0_hps_f2h_sdram0_data_waitrequest;                           // hps:f2h_sdram0_WAITREQUEST -> mm_interconnect_0:hps_f2h_sdram0_data_waitrequest
	wire   [26:0] mm_interconnect_0_hps_f2h_sdram0_data_address;                               // mm_interconnect_0:hps_f2h_sdram0_data_address -> hps:f2h_sdram0_ADDRESS
	wire          mm_interconnect_0_hps_f2h_sdram0_data_read;                                  // mm_interconnect_0:hps_f2h_sdram0_data_read -> hps:f2h_sdram0_READ
	wire   [31:0] mm_interconnect_0_hps_f2h_sdram0_data_byteenable;                            // mm_interconnect_0:hps_f2h_sdram0_data_byteenable -> hps:f2h_sdram0_BYTEENABLE
	wire          mm_interconnect_0_hps_f2h_sdram0_data_readdatavalid;                         // hps:f2h_sdram0_READDATAVALID -> mm_interconnect_0:hps_f2h_sdram0_data_readdatavalid
	wire          mm_interconnect_0_hps_f2h_sdram0_data_write;                                 // mm_interconnect_0:hps_f2h_sdram0_data_write -> hps:f2h_sdram0_WRITE
	wire  [255:0] mm_interconnect_0_hps_f2h_sdram0_data_writedata;                             // mm_interconnect_0:hps_f2h_sdram0_data_writedata -> hps:f2h_sdram0_WRITEDATA
	wire    [7:0] mm_interconnect_0_hps_f2h_sdram0_data_burstcount;                            // mm_interconnect_0:hps_f2h_sdram0_data_burstcount -> hps:f2h_sdram0_BURSTCOUNT
	wire    [1:0] hps_h2f_lw_axi_master_awburst;                                               // hps:h2f_lw_AWBURST -> mm_interconnect_1:hps_h2f_lw_axi_master_awburst
	wire    [3:0] hps_h2f_lw_axi_master_arlen;                                                 // hps:h2f_lw_ARLEN -> mm_interconnect_1:hps_h2f_lw_axi_master_arlen
	wire    [3:0] hps_h2f_lw_axi_master_wstrb;                                                 // hps:h2f_lw_WSTRB -> mm_interconnect_1:hps_h2f_lw_axi_master_wstrb
	wire          hps_h2f_lw_axi_master_wready;                                                // mm_interconnect_1:hps_h2f_lw_axi_master_wready -> hps:h2f_lw_WREADY
	wire   [11:0] hps_h2f_lw_axi_master_rid;                                                   // mm_interconnect_1:hps_h2f_lw_axi_master_rid -> hps:h2f_lw_RID
	wire          hps_h2f_lw_axi_master_rready;                                                // hps:h2f_lw_RREADY -> mm_interconnect_1:hps_h2f_lw_axi_master_rready
	wire    [3:0] hps_h2f_lw_axi_master_awlen;                                                 // hps:h2f_lw_AWLEN -> mm_interconnect_1:hps_h2f_lw_axi_master_awlen
	wire   [11:0] hps_h2f_lw_axi_master_wid;                                                   // hps:h2f_lw_WID -> mm_interconnect_1:hps_h2f_lw_axi_master_wid
	wire    [3:0] hps_h2f_lw_axi_master_arcache;                                               // hps:h2f_lw_ARCACHE -> mm_interconnect_1:hps_h2f_lw_axi_master_arcache
	wire          hps_h2f_lw_axi_master_wvalid;                                                // hps:h2f_lw_WVALID -> mm_interconnect_1:hps_h2f_lw_axi_master_wvalid
	wire   [20:0] hps_h2f_lw_axi_master_araddr;                                                // hps:h2f_lw_ARADDR -> mm_interconnect_1:hps_h2f_lw_axi_master_araddr
	wire    [2:0] hps_h2f_lw_axi_master_arprot;                                                // hps:h2f_lw_ARPROT -> mm_interconnect_1:hps_h2f_lw_axi_master_arprot
	wire    [2:0] hps_h2f_lw_axi_master_awprot;                                                // hps:h2f_lw_AWPROT -> mm_interconnect_1:hps_h2f_lw_axi_master_awprot
	wire   [31:0] hps_h2f_lw_axi_master_wdata;                                                 // hps:h2f_lw_WDATA -> mm_interconnect_1:hps_h2f_lw_axi_master_wdata
	wire          hps_h2f_lw_axi_master_arvalid;                                               // hps:h2f_lw_ARVALID -> mm_interconnect_1:hps_h2f_lw_axi_master_arvalid
	wire    [3:0] hps_h2f_lw_axi_master_awcache;                                               // hps:h2f_lw_AWCACHE -> mm_interconnect_1:hps_h2f_lw_axi_master_awcache
	wire   [11:0] hps_h2f_lw_axi_master_arid;                                                  // hps:h2f_lw_ARID -> mm_interconnect_1:hps_h2f_lw_axi_master_arid
	wire    [1:0] hps_h2f_lw_axi_master_arlock;                                                // hps:h2f_lw_ARLOCK -> mm_interconnect_1:hps_h2f_lw_axi_master_arlock
	wire    [1:0] hps_h2f_lw_axi_master_awlock;                                                // hps:h2f_lw_AWLOCK -> mm_interconnect_1:hps_h2f_lw_axi_master_awlock
	wire   [20:0] hps_h2f_lw_axi_master_awaddr;                                                // hps:h2f_lw_AWADDR -> mm_interconnect_1:hps_h2f_lw_axi_master_awaddr
	wire    [1:0] hps_h2f_lw_axi_master_bresp;                                                 // mm_interconnect_1:hps_h2f_lw_axi_master_bresp -> hps:h2f_lw_BRESP
	wire          hps_h2f_lw_axi_master_arready;                                               // mm_interconnect_1:hps_h2f_lw_axi_master_arready -> hps:h2f_lw_ARREADY
	wire   [31:0] hps_h2f_lw_axi_master_rdata;                                                 // mm_interconnect_1:hps_h2f_lw_axi_master_rdata -> hps:h2f_lw_RDATA
	wire          hps_h2f_lw_axi_master_awready;                                               // mm_interconnect_1:hps_h2f_lw_axi_master_awready -> hps:h2f_lw_AWREADY
	wire    [1:0] hps_h2f_lw_axi_master_arburst;                                               // hps:h2f_lw_ARBURST -> mm_interconnect_1:hps_h2f_lw_axi_master_arburst
	wire    [2:0] hps_h2f_lw_axi_master_arsize;                                                // hps:h2f_lw_ARSIZE -> mm_interconnect_1:hps_h2f_lw_axi_master_arsize
	wire          hps_h2f_lw_axi_master_bready;                                                // hps:h2f_lw_BREADY -> mm_interconnect_1:hps_h2f_lw_axi_master_bready
	wire          hps_h2f_lw_axi_master_rlast;                                                 // mm_interconnect_1:hps_h2f_lw_axi_master_rlast -> hps:h2f_lw_RLAST
	wire          hps_h2f_lw_axi_master_wlast;                                                 // hps:h2f_lw_WLAST -> mm_interconnect_1:hps_h2f_lw_axi_master_wlast
	wire    [1:0] hps_h2f_lw_axi_master_rresp;                                                 // mm_interconnect_1:hps_h2f_lw_axi_master_rresp -> hps:h2f_lw_RRESP
	wire   [11:0] hps_h2f_lw_axi_master_awid;                                                  // hps:h2f_lw_AWID -> mm_interconnect_1:hps_h2f_lw_axi_master_awid
	wire   [11:0] hps_h2f_lw_axi_master_bid;                                                   // mm_interconnect_1:hps_h2f_lw_axi_master_bid -> hps:h2f_lw_BID
	wire          hps_h2f_lw_axi_master_bvalid;                                                // mm_interconnect_1:hps_h2f_lw_axi_master_bvalid -> hps:h2f_lw_BVALID
	wire    [2:0] hps_h2f_lw_axi_master_awsize;                                                // hps:h2f_lw_AWSIZE -> mm_interconnect_1:hps_h2f_lw_axi_master_awsize
	wire          hps_h2f_lw_axi_master_awvalid;                                               // hps:h2f_lw_AWVALID -> mm_interconnect_1:hps_h2f_lw_axi_master_awvalid
	wire          hps_h2f_lw_axi_master_rvalid;                                                // mm_interconnect_1:hps_h2f_lw_axi_master_rvalid -> hps:h2f_lw_RVALID
	wire   [31:0] mm_interconnect_1_pipe_stage_host_ctrl_s0_readdata;                          // pipe_stage_host_ctrl:s0_readdata -> mm_interconnect_1:pipe_stage_host_ctrl_s0_readdata
	wire          mm_interconnect_1_pipe_stage_host_ctrl_s0_waitrequest;                       // pipe_stage_host_ctrl:s0_waitrequest -> mm_interconnect_1:pipe_stage_host_ctrl_s0_waitrequest
	wire          mm_interconnect_1_pipe_stage_host_ctrl_s0_debugaccess;                       // mm_interconnect_1:pipe_stage_host_ctrl_s0_debugaccess -> pipe_stage_host_ctrl:s0_debugaccess
	wire   [15:0] mm_interconnect_1_pipe_stage_host_ctrl_s0_address;                           // mm_interconnect_1:pipe_stage_host_ctrl_s0_address -> pipe_stage_host_ctrl:s0_address
	wire          mm_interconnect_1_pipe_stage_host_ctrl_s0_read;                              // mm_interconnect_1:pipe_stage_host_ctrl_s0_read -> pipe_stage_host_ctrl:s0_read
	wire    [3:0] mm_interconnect_1_pipe_stage_host_ctrl_s0_byteenable;                        // mm_interconnect_1:pipe_stage_host_ctrl_s0_byteenable -> pipe_stage_host_ctrl:s0_byteenable
	wire          mm_interconnect_1_pipe_stage_host_ctrl_s0_readdatavalid;                     // pipe_stage_host_ctrl:s0_readdatavalid -> mm_interconnect_1:pipe_stage_host_ctrl_s0_readdatavalid
	wire          mm_interconnect_1_pipe_stage_host_ctrl_s0_write;                             // mm_interconnect_1:pipe_stage_host_ctrl_s0_write -> pipe_stage_host_ctrl:s0_write
	wire   [31:0] mm_interconnect_1_pipe_stage_host_ctrl_s0_writedata;                         // mm_interconnect_1:pipe_stage_host_ctrl_s0_writedata -> pipe_stage_host_ctrl:s0_writedata
	wire    [0:0] mm_interconnect_1_pipe_stage_host_ctrl_s0_burstcount;                        // mm_interconnect_1:pipe_stage_host_ctrl_s0_burstcount -> pipe_stage_host_ctrl:s0_burstcount
	wire          pipe_stage_host_ctrl_m0_waitrequest;                                         // mm_interconnect_2:pipe_stage_host_ctrl_m0_waitrequest -> pipe_stage_host_ctrl:m0_waitrequest
	wire   [31:0] pipe_stage_host_ctrl_m0_readdata;                                            // mm_interconnect_2:pipe_stage_host_ctrl_m0_readdata -> pipe_stage_host_ctrl:m0_readdata
	wire          pipe_stage_host_ctrl_m0_debugaccess;                                         // pipe_stage_host_ctrl:m0_debugaccess -> mm_interconnect_2:pipe_stage_host_ctrl_m0_debugaccess
	wire   [15:0] pipe_stage_host_ctrl_m0_address;                                             // pipe_stage_host_ctrl:m0_address -> mm_interconnect_2:pipe_stage_host_ctrl_m0_address
	wire          pipe_stage_host_ctrl_m0_read;                                                // pipe_stage_host_ctrl:m0_read -> mm_interconnect_2:pipe_stage_host_ctrl_m0_read
	wire    [3:0] pipe_stage_host_ctrl_m0_byteenable;                                          // pipe_stage_host_ctrl:m0_byteenable -> mm_interconnect_2:pipe_stage_host_ctrl_m0_byteenable
	wire          pipe_stage_host_ctrl_m0_readdatavalid;                                       // mm_interconnect_2:pipe_stage_host_ctrl_m0_readdatavalid -> pipe_stage_host_ctrl:m0_readdatavalid
	wire   [31:0] pipe_stage_host_ctrl_m0_writedata;                                           // pipe_stage_host_ctrl:m0_writedata -> mm_interconnect_2:pipe_stage_host_ctrl_m0_writedata
	wire          pipe_stage_host_ctrl_m0_write;                                               // pipe_stage_host_ctrl:m0_write -> mm_interconnect_2:pipe_stage_host_ctrl_m0_write
	wire    [0:0] pipe_stage_host_ctrl_m0_burstcount;                                          // pipe_stage_host_ctrl:m0_burstcount -> mm_interconnect_2:pipe_stage_host_ctrl_m0_burstcount
	wire   [31:0] mm_interconnect_2_acl_kernel_interface_ctrl_readdata;                        // acl_kernel_interface:ctrl_readdata -> mm_interconnect_2:acl_kernel_interface_ctrl_readdata
	wire          mm_interconnect_2_acl_kernel_interface_ctrl_waitrequest;                     // acl_kernel_interface:ctrl_waitrequest -> mm_interconnect_2:acl_kernel_interface_ctrl_waitrequest
	wire          mm_interconnect_2_acl_kernel_interface_ctrl_debugaccess;                     // mm_interconnect_2:acl_kernel_interface_ctrl_debugaccess -> acl_kernel_interface:ctrl_debugaccess
	wire   [13:0] mm_interconnect_2_acl_kernel_interface_ctrl_address;                         // mm_interconnect_2:acl_kernel_interface_ctrl_address -> acl_kernel_interface:ctrl_address
	wire          mm_interconnect_2_acl_kernel_interface_ctrl_read;                            // mm_interconnect_2:acl_kernel_interface_ctrl_read -> acl_kernel_interface:ctrl_read
	wire    [3:0] mm_interconnect_2_acl_kernel_interface_ctrl_byteenable;                      // mm_interconnect_2:acl_kernel_interface_ctrl_byteenable -> acl_kernel_interface:ctrl_byteenable
	wire          mm_interconnect_2_acl_kernel_interface_ctrl_readdatavalid;                   // acl_kernel_interface:ctrl_readdatavalid -> mm_interconnect_2:acl_kernel_interface_ctrl_readdatavalid
	wire          mm_interconnect_2_acl_kernel_interface_ctrl_write;                           // mm_interconnect_2:acl_kernel_interface_ctrl_write -> acl_kernel_interface:ctrl_write
	wire   [31:0] mm_interconnect_2_acl_kernel_interface_ctrl_writedata;                       // mm_interconnect_2:acl_kernel_interface_ctrl_writedata -> acl_kernel_interface:ctrl_writedata
	wire    [0:0] mm_interconnect_2_acl_kernel_interface_ctrl_burstcount;                      // mm_interconnect_2:acl_kernel_interface_ctrl_burstcount -> acl_kernel_interface:ctrl_burstcount
	wire   [31:0] mm_interconnect_2_version_id_s_readdata;                                     // version_id:slave_readdata -> mm_interconnect_2:version_id_s_readdata
	wire          mm_interconnect_2_version_id_s_read;                                         // mm_interconnect_2:version_id_s_read -> version_id:slave_read
	wire          clock_cross_kernel_mem1_m0_waitrequest;                                      // mm_interconnect_3:clock_cross_kernel_mem1_m0_waitrequest -> clock_cross_kernel_mem1:m0_waitrequest
	wire  [255:0] clock_cross_kernel_mem1_m0_readdata;                                         // mm_interconnect_3:clock_cross_kernel_mem1_m0_readdata -> clock_cross_kernel_mem1:m0_readdata
	wire          clock_cross_kernel_mem1_m0_debugaccess;                                      // clock_cross_kernel_mem1:m0_debugaccess -> mm_interconnect_3:clock_cross_kernel_mem1_m0_debugaccess
	wire   [24:0] clock_cross_kernel_mem1_m0_address;                                          // clock_cross_kernel_mem1:m0_address -> mm_interconnect_3:clock_cross_kernel_mem1_m0_address
	wire          clock_cross_kernel_mem1_m0_read;                                             // clock_cross_kernel_mem1:m0_read -> mm_interconnect_3:clock_cross_kernel_mem1_m0_read
	wire   [31:0] clock_cross_kernel_mem1_m0_byteenable;                                       // clock_cross_kernel_mem1:m0_byteenable -> mm_interconnect_3:clock_cross_kernel_mem1_m0_byteenable
	wire          clock_cross_kernel_mem1_m0_readdatavalid;                                    // mm_interconnect_3:clock_cross_kernel_mem1_m0_readdatavalid -> clock_cross_kernel_mem1:m0_readdatavalid
	wire  [255:0] clock_cross_kernel_mem1_m0_writedata;                                        // clock_cross_kernel_mem1:m0_writedata -> mm_interconnect_3:clock_cross_kernel_mem1_m0_writedata
	wire          clock_cross_kernel_mem1_m0_write;                                            // clock_cross_kernel_mem1:m0_write -> mm_interconnect_3:clock_cross_kernel_mem1_m0_write
	wire    [4:0] clock_cross_kernel_mem1_m0_burstcount;                                       // clock_cross_kernel_mem1:m0_burstcount -> mm_interconnect_3:clock_cross_kernel_mem1_m0_burstcount
	wire  [255:0] mm_interconnect_3_address_span_extender_kernel_windowed_slave_readdata;      // address_span_extender_kernel:avs_s0_readdata -> mm_interconnect_3:address_span_extender_kernel_windowed_slave_readdata
	wire          mm_interconnect_3_address_span_extender_kernel_windowed_slave_waitrequest;   // address_span_extender_kernel:avs_s0_waitrequest -> mm_interconnect_3:address_span_extender_kernel_windowed_slave_waitrequest
	wire   [24:0] mm_interconnect_3_address_span_extender_kernel_windowed_slave_address;       // mm_interconnect_3:address_span_extender_kernel_windowed_slave_address -> address_span_extender_kernel:avs_s0_address
	wire          mm_interconnect_3_address_span_extender_kernel_windowed_slave_read;          // mm_interconnect_3:address_span_extender_kernel_windowed_slave_read -> address_span_extender_kernel:avs_s0_read
	wire   [31:0] mm_interconnect_3_address_span_extender_kernel_windowed_slave_byteenable;    // mm_interconnect_3:address_span_extender_kernel_windowed_slave_byteenable -> address_span_extender_kernel:avs_s0_byteenable
	wire          mm_interconnect_3_address_span_extender_kernel_windowed_slave_readdatavalid; // address_span_extender_kernel:avs_s0_readdatavalid -> mm_interconnect_3:address_span_extender_kernel_windowed_slave_readdatavalid
	wire          mm_interconnect_3_address_span_extender_kernel_windowed_slave_write;         // mm_interconnect_3:address_span_extender_kernel_windowed_slave_write -> address_span_extender_kernel:avs_s0_write
	wire  [255:0] mm_interconnect_3_address_span_extender_kernel_windowed_slave_writedata;     // mm_interconnect_3:address_span_extender_kernel_windowed_slave_writedata -> address_span_extender_kernel:avs_s0_writedata
	wire    [4:0] mm_interconnect_3_address_span_extender_kernel_windowed_slave_burstcount;    // mm_interconnect_3:address_span_extender_kernel_windowed_slave_burstcount -> address_span_extender_kernel:avs_s0_burstcount
	wire          irq_mapper_receiver0_irq;                                                    // acl_kernel_interface:kernel_irq_to_host_irq -> irq_mapper:receiver0_irq
	wire   [31:0] hps_f2h_irq0_irq;                                                            // irq_mapper:sender_irq -> hps:f2h_irq_p0
	wire   [31:0] hps_f2h_irq1_irq;                                                            // irq_mapper_001:sender_irq -> hps:f2h_irq_p1
	wire          rst_controller_reset_out_reset;                                              // rst_controller:reset_out -> [acl_kernel_clk:reset_reset_n, acl_kernel_interface:reset_reset_n, acl_kernel_interface:sw_reset_in_reset, mm_interconnect_1:pipe_stage_host_ctrl_reset_reset_bridge_in_reset_reset, mm_interconnect_2:pipe_stage_host_ctrl_reset_reset_bridge_in_reset_reset, pipe_stage_host_ctrl:reset, version_id:resetn]
	wire          rst_controller_001_reset_out_reset;                                          // rst_controller_001:reset_out -> [address_span_extender_kernel:reset, clock_cross_kernel_mem1:m0_reset, mm_interconnect_0:address_span_extender_kernel_reset_reset_bridge_in_reset_reset, mm_interconnect_3:clock_cross_kernel_mem1_m0_reset_reset_bridge_in_reset_reset]
	wire          acl_kernel_interface_sw_reset_export_reset;                                  // acl_kernel_interface:sw_reset_export_reset_n -> rst_controller_001:reset_in0
	wire          rst_controller_002_reset_out_reset;                                          // rst_controller_002:reset_out -> mm_interconnect_0:hps_f2h_sdram0_data_translator_reset_reset_bridge_in_reset_reset
	wire          hps_h2f_reset_reset;                                                         // hps:h2f_rst_n -> [rst_controller_002:reset_in0, rst_controller_003:reset_in0]
	wire          rst_controller_003_reset_out_reset;                                          // rst_controller_003:reset_out -> mm_interconnect_1:hps_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset

	system_acl_iface_acl_kernel_clk acl_kernel_clk (
		.pll_refclk_clk           (kernel_pll_refclk_clk),                   //        pll_refclk.clk
		.clk_clk                  (config_clk_clk),                          //               clk.clk
		.reset_reset_n            (~rst_controller_reset_out_reset),         //             reset.reset_n
		.ctrl_waitrequest         (),                                        //              ctrl.waitrequest
		.ctrl_readdata            (),                                        //                  .readdata
		.ctrl_readdatavalid       (),                                        //                  .readdatavalid
		.ctrl_burstcount          (),                                        //                  .burstcount
		.ctrl_writedata           (),                                        //                  .writedata
		.ctrl_address             (),                                        //                  .address
		.ctrl_write               (),                                        //                  .write
		.ctrl_read                (),                                        //                  .read
		.ctrl_byteenable          (),                                        //                  .byteenable
		.ctrl_debugaccess         (),                                        //                  .debugaccess
		.kernel_clk_clk           (kernel_clk_clk),                          //        kernel_clk.clk
		.kernel_clk2x_clk         (kernel_clk2x_clk),                        //      kernel_clk2x.clk
		.kernel_pll_locked_export (acl_kernel_clk_kernel_pll_locked_export)  // kernel_pll_locked.export
	);

	system_acl_iface_acl_kernel_interface acl_kernel_interface (
		.clk_clk                       (config_clk_clk),                                            //                      clk.clk
		.reset_reset_n                 (~rst_controller_reset_out_reset),                           //                    reset.reset_n
		.ctrl_waitrequest              (mm_interconnect_2_acl_kernel_interface_ctrl_waitrequest),   //                     ctrl.waitrequest
		.ctrl_readdata                 (mm_interconnect_2_acl_kernel_interface_ctrl_readdata),      //                         .readdata
		.ctrl_readdatavalid            (mm_interconnect_2_acl_kernel_interface_ctrl_readdatavalid), //                         .readdatavalid
		.ctrl_burstcount               (mm_interconnect_2_acl_kernel_interface_ctrl_burstcount),    //                         .burstcount
		.ctrl_writedata                (mm_interconnect_2_acl_kernel_interface_ctrl_writedata),     //                         .writedata
		.ctrl_address                  (mm_interconnect_2_acl_kernel_interface_ctrl_address),       //                         .address
		.ctrl_write                    (mm_interconnect_2_acl_kernel_interface_ctrl_write),         //                         .write
		.ctrl_read                     (mm_interconnect_2_acl_kernel_interface_ctrl_read),          //                         .read
		.ctrl_byteenable               (mm_interconnect_2_acl_kernel_interface_ctrl_byteenable),    //                         .byteenable
		.ctrl_debugaccess              (mm_interconnect_2_acl_kernel_interface_ctrl_debugaccess),   //                         .debugaccess
		.kernel_cra_waitrequest        (kernel_cra_waitrequest),                                    //               kernel_cra.waitrequest
		.kernel_cra_readdata           (kernel_cra_readdata),                                       //                         .readdata
		.kernel_cra_readdatavalid      (kernel_cra_readdatavalid),                                  //                         .readdatavalid
		.kernel_cra_burstcount         (kernel_cra_burstcount),                                     //                         .burstcount
		.kernel_cra_writedata          (kernel_cra_writedata),                                      //                         .writedata
		.kernel_cra_address            (kernel_cra_address),                                        //                         .address
		.kernel_cra_write              (kernel_cra_write),                                          //                         .write
		.kernel_cra_read               (kernel_cra_read),                                           //                         .read
		.kernel_cra_byteenable         (kernel_cra_byteenable),                                     //                         .byteenable
		.kernel_cra_debugaccess        (kernel_cra_debugaccess),                                    //                         .debugaccess
		.kernel_irq_from_kernel_irq    (kernel_irq_irq),                                            //   kernel_irq_from_kernel.irq
		.acl_bsp_memorg_kernel_mode    (acl_internal_memorg_kernel_mode),                           //    acl_bsp_memorg_kernel.mode
		.acl_bsp_memorg_host0x018_mode (),                                                          // acl_bsp_memorg_host0x018.mode
		.sw_reset_in_reset             (rst_controller_reset_out_reset),                            //              sw_reset_in.reset
		.kernel_clk_clk                (kernel_clk_clk),                                            //               kernel_clk.clk
		.sw_reset_export_reset_n       (acl_kernel_interface_sw_reset_export_reset),                //          sw_reset_export.reset_n
		.kernel_reset_reset_n          (kernel_reset_reset_n),                                      //             kernel_reset.reset_n
		.kernel_irq_to_host_irq        (irq_mapper_receiver0_irq)                                   //       kernel_irq_to_host.irq
	);

	altera_address_span_extender #(
		.DATA_WIDTH           (256),
		.BYTEENABLE_WIDTH     (32),
		.MASTER_ADDRESS_WIDTH (32),
		.SLAVE_ADDRESS_WIDTH  (25),
		.SLAVE_ADDRESS_SHIFT  (5),
		.BURSTCOUNT_WIDTH     (5),
		.CNTL_ADDRESS_WIDTH   (1),
		.SUB_WINDOW_COUNT     (1),
		.MASTER_ADDRESS_DEF   (64'b0000000000000000000000000000000000000000000000000000000000000000)
	) address_span_extender_kernel (
		.clk                  (pll_outclk0_clk),                                                             //           clock.clk
		.reset                (rst_controller_001_reset_out_reset),                                          //           reset.reset
		.avs_s0_address       (mm_interconnect_3_address_span_extender_kernel_windowed_slave_address),       //  windowed_slave.address
		.avs_s0_read          (mm_interconnect_3_address_span_extender_kernel_windowed_slave_read),          //                .read
		.avs_s0_readdata      (mm_interconnect_3_address_span_extender_kernel_windowed_slave_readdata),      //                .readdata
		.avs_s0_write         (mm_interconnect_3_address_span_extender_kernel_windowed_slave_write),         //                .write
		.avs_s0_writedata     (mm_interconnect_3_address_span_extender_kernel_windowed_slave_writedata),     //                .writedata
		.avs_s0_readdatavalid (mm_interconnect_3_address_span_extender_kernel_windowed_slave_readdatavalid), //                .readdatavalid
		.avs_s0_waitrequest   (mm_interconnect_3_address_span_extender_kernel_windowed_slave_waitrequest),   //                .waitrequest
		.avs_s0_byteenable    (mm_interconnect_3_address_span_extender_kernel_windowed_slave_byteenable),    //                .byteenable
		.avs_s0_burstcount    (mm_interconnect_3_address_span_extender_kernel_windowed_slave_burstcount),    //                .burstcount
		.avm_m0_address       (address_span_extender_kernel_expanded_master_address),                        // expanded_master.address
		.avm_m0_read          (address_span_extender_kernel_expanded_master_read),                           //                .read
		.avm_m0_waitrequest   (address_span_extender_kernel_expanded_master_waitrequest),                    //                .waitrequest
		.avm_m0_readdata      (address_span_extender_kernel_expanded_master_readdata),                       //                .readdata
		.avm_m0_write         (address_span_extender_kernel_expanded_master_write),                          //                .write
		.avm_m0_writedata     (address_span_extender_kernel_expanded_master_writedata),                      //                .writedata
		.avm_m0_readdatavalid (address_span_extender_kernel_expanded_master_readdatavalid),                  //                .readdatavalid
		.avm_m0_byteenable    (address_span_extender_kernel_expanded_master_byteenable),                     //                .byteenable
		.avm_m0_burstcount    (address_span_extender_kernel_expanded_master_burstcount),                     //                .burstcount
		.avs_cntl_address     (1'b0),                                                                        //     (terminated)
		.avs_cntl_read        (1'b0),                                                                        //     (terminated)
		.avs_cntl_readdata    (),                                                                            //     (terminated)
		.avs_cntl_write       (1'b0),                                                                        //     (terminated)
		.avs_cntl_writedata   (64'b0000000000000000000000000000000000000000000000000000000000000000),        //     (terminated)
		.avs_cntl_byteenable  (8'b00000000)                                                                  //     (terminated)
	);

	altera_avalon_mm_clock_crossing_bridge #(
		.DATA_WIDTH          (256),
		.SYMBOL_WIDTH        (8),
		.HDL_ADDR_WIDTH      (25),
		.BURSTCOUNT_WIDTH    (5),
		.COMMAND_FIFO_DEPTH  (64),
		.RESPONSE_FIFO_DEPTH (64),
		.MASTER_SYNC_DEPTH   (2),
		.SLAVE_SYNC_DEPTH    (2)
	) clock_cross_kernel_mem1 (
		.m0_clk           (pll_outclk0_clk),                          //   m0_clk.clk
		.m0_reset         (rst_controller_001_reset_out_reset),       // m0_reset.reset
		.s0_clk           (kernel_clk_clk),                           //   s0_clk.clk
		.s0_reset         (~kernel_reset_reset_n),                    // s0_reset.reset
		.s0_waitrequest   (kernel_mem0_waitrequest),                  //       s0.waitrequest
		.s0_readdata      (kernel_mem0_readdata),                     //         .readdata
		.s0_readdatavalid (kernel_mem0_readdatavalid),                //         .readdatavalid
		.s0_burstcount    (kernel_mem0_burstcount),                   //         .burstcount
		.s0_writedata     (kernel_mem0_writedata),                    //         .writedata
		.s0_address       (kernel_mem0_address),                      //         .address
		.s0_write         (kernel_mem0_write),                        //         .write
		.s0_read          (kernel_mem0_read),                         //         .read
		.s0_byteenable    (kernel_mem0_byteenable),                   //         .byteenable
		.s0_debugaccess   (kernel_mem0_debugaccess),                  //         .debugaccess
		.m0_waitrequest   (clock_cross_kernel_mem1_m0_waitrequest),   //       m0.waitrequest
		.m0_readdata      (clock_cross_kernel_mem1_m0_readdata),      //         .readdata
		.m0_readdatavalid (clock_cross_kernel_mem1_m0_readdatavalid), //         .readdatavalid
		.m0_burstcount    (clock_cross_kernel_mem1_m0_burstcount),    //         .burstcount
		.m0_writedata     (clock_cross_kernel_mem1_m0_writedata),     //         .writedata
		.m0_address       (clock_cross_kernel_mem1_m0_address),       //         .address
		.m0_write         (clock_cross_kernel_mem1_m0_write),         //         .write
		.m0_read          (clock_cross_kernel_mem1_m0_read),          //         .read
		.m0_byteenable    (clock_cross_kernel_mem1_m0_byteenable),    //         .byteenable
		.m0_debugaccess   (clock_cross_kernel_mem1_m0_debugaccess)    //         .debugaccess
	);

	system_acl_iface_hps #(
		.F2S_Width (0),
		.S2F_Width (0)
	) hps (
		.mem_a                    (memory_mem_a),                                        //            memory.mem_a
		.mem_ba                   (memory_mem_ba),                                       //                  .mem_ba
		.mem_ck                   (memory_mem_ck),                                       //                  .mem_ck
		.mem_ck_n                 (memory_mem_ck_n),                                     //                  .mem_ck_n
		.mem_cke                  (memory_mem_cke),                                      //                  .mem_cke
		.mem_cs_n                 (memory_mem_cs_n),                                     //                  .mem_cs_n
		.mem_ras_n                (memory_mem_ras_n),                                    //                  .mem_ras_n
		.mem_cas_n                (memory_mem_cas_n),                                    //                  .mem_cas_n
		.mem_we_n                 (memory_mem_we_n),                                     //                  .mem_we_n
		.mem_reset_n              (memory_mem_reset_n),                                  //                  .mem_reset_n
		.mem_dq                   (memory_mem_dq),                                       //                  .mem_dq
		.mem_dqs                  (memory_mem_dqs),                                      //                  .mem_dqs
		.mem_dqs_n                (memory_mem_dqs_n),                                    //                  .mem_dqs_n
		.mem_odt                  (memory_mem_odt),                                      //                  .mem_odt
		.mem_dm                   (memory_mem_dm),                                       //                  .mem_dm
		.oct_rzqin                (memory_oct_rzqin),                                    //                  .oct_rzqin
		.hps_io_emac1_inst_TX_CLK (peripheral_hps_io_emac1_inst_TX_CLK),                 //            hps_io.hps_io_emac1_inst_TX_CLK
		.hps_io_emac1_inst_TXD0   (peripheral_hps_io_emac1_inst_TXD0),                   //                  .hps_io_emac1_inst_TXD0
		.hps_io_emac1_inst_TXD1   (peripheral_hps_io_emac1_inst_TXD1),                   //                  .hps_io_emac1_inst_TXD1
		.hps_io_emac1_inst_TXD2   (peripheral_hps_io_emac1_inst_TXD2),                   //                  .hps_io_emac1_inst_TXD2
		.hps_io_emac1_inst_TXD3   (peripheral_hps_io_emac1_inst_TXD3),                   //                  .hps_io_emac1_inst_TXD3
		.hps_io_emac1_inst_RXD0   (peripheral_hps_io_emac1_inst_RXD0),                   //                  .hps_io_emac1_inst_RXD0
		.hps_io_emac1_inst_MDIO   (peripheral_hps_io_emac1_inst_MDIO),                   //                  .hps_io_emac1_inst_MDIO
		.hps_io_emac1_inst_MDC    (peripheral_hps_io_emac1_inst_MDC),                    //                  .hps_io_emac1_inst_MDC
		.hps_io_emac1_inst_RX_CTL (peripheral_hps_io_emac1_inst_RX_CTL),                 //                  .hps_io_emac1_inst_RX_CTL
		.hps_io_emac1_inst_TX_CTL (peripheral_hps_io_emac1_inst_TX_CTL),                 //                  .hps_io_emac1_inst_TX_CTL
		.hps_io_emac1_inst_RX_CLK (peripheral_hps_io_emac1_inst_RX_CLK),                 //                  .hps_io_emac1_inst_RX_CLK
		.hps_io_emac1_inst_RXD1   (peripheral_hps_io_emac1_inst_RXD1),                   //                  .hps_io_emac1_inst_RXD1
		.hps_io_emac1_inst_RXD2   (peripheral_hps_io_emac1_inst_RXD2),                   //                  .hps_io_emac1_inst_RXD2
		.hps_io_emac1_inst_RXD3   (peripheral_hps_io_emac1_inst_RXD3),                   //                  .hps_io_emac1_inst_RXD3
		.hps_io_sdio_inst_CMD     (peripheral_hps_io_sdio_inst_CMD),                     //                  .hps_io_sdio_inst_CMD
		.hps_io_sdio_inst_D0      (peripheral_hps_io_sdio_inst_D0),                      //                  .hps_io_sdio_inst_D0
		.hps_io_sdio_inst_D1      (peripheral_hps_io_sdio_inst_D1),                      //                  .hps_io_sdio_inst_D1
		.hps_io_sdio_inst_CLK     (peripheral_hps_io_sdio_inst_CLK),                     //                  .hps_io_sdio_inst_CLK
		.hps_io_sdio_inst_D2      (peripheral_hps_io_sdio_inst_D2),                      //                  .hps_io_sdio_inst_D2
		.hps_io_sdio_inst_D3      (peripheral_hps_io_sdio_inst_D3),                      //                  .hps_io_sdio_inst_D3
		.hps_io_usb1_inst_D0      (peripheral_hps_io_usb1_inst_D0),                      //                  .hps_io_usb1_inst_D0
		.hps_io_usb1_inst_D1      (peripheral_hps_io_usb1_inst_D1),                      //                  .hps_io_usb1_inst_D1
		.hps_io_usb1_inst_D2      (peripheral_hps_io_usb1_inst_D2),                      //                  .hps_io_usb1_inst_D2
		.hps_io_usb1_inst_D3      (peripheral_hps_io_usb1_inst_D3),                      //                  .hps_io_usb1_inst_D3
		.hps_io_usb1_inst_D4      (peripheral_hps_io_usb1_inst_D4),                      //                  .hps_io_usb1_inst_D4
		.hps_io_usb1_inst_D5      (peripheral_hps_io_usb1_inst_D5),                      //                  .hps_io_usb1_inst_D5
		.hps_io_usb1_inst_D6      (peripheral_hps_io_usb1_inst_D6),                      //                  .hps_io_usb1_inst_D6
		.hps_io_usb1_inst_D7      (peripheral_hps_io_usb1_inst_D7),                      //                  .hps_io_usb1_inst_D7
		.hps_io_usb1_inst_CLK     (peripheral_hps_io_usb1_inst_CLK),                     //                  .hps_io_usb1_inst_CLK
		.hps_io_usb1_inst_STP     (peripheral_hps_io_usb1_inst_STP),                     //                  .hps_io_usb1_inst_STP
		.hps_io_usb1_inst_DIR     (peripheral_hps_io_usb1_inst_DIR),                     //                  .hps_io_usb1_inst_DIR
		.hps_io_usb1_inst_NXT     (peripheral_hps_io_usb1_inst_NXT),                     //                  .hps_io_usb1_inst_NXT
		.hps_io_uart0_inst_RX     (peripheral_hps_io_uart0_inst_RX),                     //                  .hps_io_uart0_inst_RX
		.hps_io_uart0_inst_TX     (peripheral_hps_io_uart0_inst_TX),                     //                  .hps_io_uart0_inst_TX
		.hps_io_i2c1_inst_SDA     (peripheral_hps_io_i2c1_inst_SDA),                     //                  .hps_io_i2c1_inst_SDA
		.hps_io_i2c1_inst_SCL     (peripheral_hps_io_i2c1_inst_SCL),                     //                  .hps_io_i2c1_inst_SCL
		.hps_io_gpio_inst_GPIO53  (peripheral_hps_io_gpio_inst_GPIO53),                  //                  .hps_io_gpio_inst_GPIO53
		.h2f_rst_n                (hps_h2f_reset_reset),                                 //         h2f_reset.reset_n
		.f2h_sdram0_clk           (pll_outclk0_clk),                                     //  f2h_sdram0_clock.clk
		.f2h_sdram0_ADDRESS       (mm_interconnect_0_hps_f2h_sdram0_data_address),       //   f2h_sdram0_data.address
		.f2h_sdram0_BURSTCOUNT    (mm_interconnect_0_hps_f2h_sdram0_data_burstcount),    //                  .burstcount
		.f2h_sdram0_WAITREQUEST   (mm_interconnect_0_hps_f2h_sdram0_data_waitrequest),   //                  .waitrequest
		.f2h_sdram0_READDATA      (mm_interconnect_0_hps_f2h_sdram0_data_readdata),      //                  .readdata
		.f2h_sdram0_READDATAVALID (mm_interconnect_0_hps_f2h_sdram0_data_readdatavalid), //                  .readdatavalid
		.f2h_sdram0_READ          (mm_interconnect_0_hps_f2h_sdram0_data_read),          //                  .read
		.f2h_sdram0_WRITEDATA     (mm_interconnect_0_hps_f2h_sdram0_data_writedata),     //                  .writedata
		.f2h_sdram0_BYTEENABLE    (mm_interconnect_0_hps_f2h_sdram0_data_byteenable),    //                  .byteenable
		.f2h_sdram0_WRITE         (mm_interconnect_0_hps_f2h_sdram0_data_write),         //                  .write
		.h2f_lw_axi_clk           (config_clk_clk),                                      //  h2f_lw_axi_clock.clk
		.h2f_lw_AWID              (hps_h2f_lw_axi_master_awid),                          // h2f_lw_axi_master.awid
		.h2f_lw_AWADDR            (hps_h2f_lw_axi_master_awaddr),                        //                  .awaddr
		.h2f_lw_AWLEN             (hps_h2f_lw_axi_master_awlen),                         //                  .awlen
		.h2f_lw_AWSIZE            (hps_h2f_lw_axi_master_awsize),                        //                  .awsize
		.h2f_lw_AWBURST           (hps_h2f_lw_axi_master_awburst),                       //                  .awburst
		.h2f_lw_AWLOCK            (hps_h2f_lw_axi_master_awlock),                        //                  .awlock
		.h2f_lw_AWCACHE           (hps_h2f_lw_axi_master_awcache),                       //                  .awcache
		.h2f_lw_AWPROT            (hps_h2f_lw_axi_master_awprot),                        //                  .awprot
		.h2f_lw_AWVALID           (hps_h2f_lw_axi_master_awvalid),                       //                  .awvalid
		.h2f_lw_AWREADY           (hps_h2f_lw_axi_master_awready),                       //                  .awready
		.h2f_lw_WID               (hps_h2f_lw_axi_master_wid),                           //                  .wid
		.h2f_lw_WDATA             (hps_h2f_lw_axi_master_wdata),                         //                  .wdata
		.h2f_lw_WSTRB             (hps_h2f_lw_axi_master_wstrb),                         //                  .wstrb
		.h2f_lw_WLAST             (hps_h2f_lw_axi_master_wlast),                         //                  .wlast
		.h2f_lw_WVALID            (hps_h2f_lw_axi_master_wvalid),                        //                  .wvalid
		.h2f_lw_WREADY            (hps_h2f_lw_axi_master_wready),                        //                  .wready
		.h2f_lw_BID               (hps_h2f_lw_axi_master_bid),                           //                  .bid
		.h2f_lw_BRESP             (hps_h2f_lw_axi_master_bresp),                         //                  .bresp
		.h2f_lw_BVALID            (hps_h2f_lw_axi_master_bvalid),                        //                  .bvalid
		.h2f_lw_BREADY            (hps_h2f_lw_axi_master_bready),                        //                  .bready
		.h2f_lw_ARID              (hps_h2f_lw_axi_master_arid),                          //                  .arid
		.h2f_lw_ARADDR            (hps_h2f_lw_axi_master_araddr),                        //                  .araddr
		.h2f_lw_ARLEN             (hps_h2f_lw_axi_master_arlen),                         //                  .arlen
		.h2f_lw_ARSIZE            (hps_h2f_lw_axi_master_arsize),                        //                  .arsize
		.h2f_lw_ARBURST           (hps_h2f_lw_axi_master_arburst),                       //                  .arburst
		.h2f_lw_ARLOCK            (hps_h2f_lw_axi_master_arlock),                        //                  .arlock
		.h2f_lw_ARCACHE           (hps_h2f_lw_axi_master_arcache),                       //                  .arcache
		.h2f_lw_ARPROT            (hps_h2f_lw_axi_master_arprot),                        //                  .arprot
		.h2f_lw_ARVALID           (hps_h2f_lw_axi_master_arvalid),                       //                  .arvalid
		.h2f_lw_ARREADY           (hps_h2f_lw_axi_master_arready),                       //                  .arready
		.h2f_lw_RID               (hps_h2f_lw_axi_master_rid),                           //                  .rid
		.h2f_lw_RDATA             (hps_h2f_lw_axi_master_rdata),                         //                  .rdata
		.h2f_lw_RRESP             (hps_h2f_lw_axi_master_rresp),                         //                  .rresp
		.h2f_lw_RLAST             (hps_h2f_lw_axi_master_rlast),                         //                  .rlast
		.h2f_lw_RVALID            (hps_h2f_lw_axi_master_rvalid),                        //                  .rvalid
		.h2f_lw_RREADY            (hps_h2f_lw_axi_master_rready),                        //                  .rready
		.f2h_irq_p0               (hps_f2h_irq0_irq),                                    //          f2h_irq0.irq
		.f2h_irq_p1               (hps_f2h_irq1_irq)                                     //          f2h_irq1.irq
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (32),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (16),
		.BURSTCOUNT_WIDTH  (1),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) pipe_stage_host_ctrl (
		.clk              (config_clk_clk),                                          //   clk.clk
		.reset            (rst_controller_reset_out_reset),                          // reset.reset
		.s0_waitrequest   (mm_interconnect_1_pipe_stage_host_ctrl_s0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (mm_interconnect_1_pipe_stage_host_ctrl_s0_readdata),      //      .readdata
		.s0_readdatavalid (mm_interconnect_1_pipe_stage_host_ctrl_s0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (mm_interconnect_1_pipe_stage_host_ctrl_s0_burstcount),    //      .burstcount
		.s0_writedata     (mm_interconnect_1_pipe_stage_host_ctrl_s0_writedata),     //      .writedata
		.s0_address       (mm_interconnect_1_pipe_stage_host_ctrl_s0_address),       //      .address
		.s0_write         (mm_interconnect_1_pipe_stage_host_ctrl_s0_write),         //      .write
		.s0_read          (mm_interconnect_1_pipe_stage_host_ctrl_s0_read),          //      .read
		.s0_byteenable    (mm_interconnect_1_pipe_stage_host_ctrl_s0_byteenable),    //      .byteenable
		.s0_debugaccess   (mm_interconnect_1_pipe_stage_host_ctrl_s0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (pipe_stage_host_ctrl_m0_waitrequest),                     //    m0.waitrequest
		.m0_readdata      (pipe_stage_host_ctrl_m0_readdata),                        //      .readdata
		.m0_readdatavalid (pipe_stage_host_ctrl_m0_readdatavalid),                   //      .readdatavalid
		.m0_burstcount    (pipe_stage_host_ctrl_m0_burstcount),                      //      .burstcount
		.m0_writedata     (pipe_stage_host_ctrl_m0_writedata),                       //      .writedata
		.m0_address       (pipe_stage_host_ctrl_m0_address),                         //      .address
		.m0_write         (pipe_stage_host_ctrl_m0_write),                           //      .write
		.m0_read          (pipe_stage_host_ctrl_m0_read),                            //      .read
		.m0_byteenable    (pipe_stage_host_ctrl_m0_byteenable),                      //      .byteenable
		.m0_debugaccess   (pipe_stage_host_ctrl_m0_debugaccess),                     //      .debugaccess
		.s0_response      (),                                                        // (terminated)
		.m0_response      (2'b00)                                                    // (terminated)
	);

	system_acl_iface_pll pll (
		.refclk   (config_clk_clk),  //  refclk.clk
		.rst      (~reset_n),        //   reset.reset
		.outclk_0 (pll_outclk0_clk), // outclk0.clk
		.locked   ()                 // (terminated)
	);

	version_id #(
		.WIDTH      (32),
		.VERSION_ID (-1597521440)
	) version_id (
		.clk            (config_clk_clk),                          //       clk.clk
		.resetn         (~rst_controller_reset_out_reset),         // clk_reset.reset_n
		.slave_read     (mm_interconnect_2_version_id_s_read),     //         s.read
		.slave_readdata (mm_interconnect_2_version_id_s_readdata)  //          .readdata
	);

	system_acl_iface_mm_interconnect_0 mm_interconnect_0 (
		.pll_outclk0_clk                                                  (pll_outclk0_clk),                                            //                                                pll_outclk0.clk
		.address_span_extender_kernel_reset_reset_bridge_in_reset_reset   (rst_controller_001_reset_out_reset),                         //   address_span_extender_kernel_reset_reset_bridge_in_reset.reset
		.hps_f2h_sdram0_data_translator_reset_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),                         // hps_f2h_sdram0_data_translator_reset_reset_bridge_in_reset.reset
		.address_span_extender_kernel_expanded_master_address             (address_span_extender_kernel_expanded_master_address),       //               address_span_extender_kernel_expanded_master.address
		.address_span_extender_kernel_expanded_master_waitrequest         (address_span_extender_kernel_expanded_master_waitrequest),   //                                                           .waitrequest
		.address_span_extender_kernel_expanded_master_burstcount          (address_span_extender_kernel_expanded_master_burstcount),    //                                                           .burstcount
		.address_span_extender_kernel_expanded_master_byteenable          (address_span_extender_kernel_expanded_master_byteenable),    //                                                           .byteenable
		.address_span_extender_kernel_expanded_master_read                (address_span_extender_kernel_expanded_master_read),          //                                                           .read
		.address_span_extender_kernel_expanded_master_readdata            (address_span_extender_kernel_expanded_master_readdata),      //                                                           .readdata
		.address_span_extender_kernel_expanded_master_readdatavalid       (address_span_extender_kernel_expanded_master_readdatavalid), //                                                           .readdatavalid
		.address_span_extender_kernel_expanded_master_write               (address_span_extender_kernel_expanded_master_write),         //                                                           .write
		.address_span_extender_kernel_expanded_master_writedata           (address_span_extender_kernel_expanded_master_writedata),     //                                                           .writedata
		.hps_f2h_sdram0_data_address                                      (mm_interconnect_0_hps_f2h_sdram0_data_address),              //                                        hps_f2h_sdram0_data.address
		.hps_f2h_sdram0_data_write                                        (mm_interconnect_0_hps_f2h_sdram0_data_write),                //                                                           .write
		.hps_f2h_sdram0_data_read                                         (mm_interconnect_0_hps_f2h_sdram0_data_read),                 //                                                           .read
		.hps_f2h_sdram0_data_readdata                                     (mm_interconnect_0_hps_f2h_sdram0_data_readdata),             //                                                           .readdata
		.hps_f2h_sdram0_data_writedata                                    (mm_interconnect_0_hps_f2h_sdram0_data_writedata),            //                                                           .writedata
		.hps_f2h_sdram0_data_burstcount                                   (mm_interconnect_0_hps_f2h_sdram0_data_burstcount),           //                                                           .burstcount
		.hps_f2h_sdram0_data_byteenable                                   (mm_interconnect_0_hps_f2h_sdram0_data_byteenable),           //                                                           .byteenable
		.hps_f2h_sdram0_data_readdatavalid                                (mm_interconnect_0_hps_f2h_sdram0_data_readdatavalid),        //                                                           .readdatavalid
		.hps_f2h_sdram0_data_waitrequest                                  (mm_interconnect_0_hps_f2h_sdram0_data_waitrequest)           //                                                           .waitrequest
	);

	system_acl_iface_mm_interconnect_1 mm_interconnect_1 (
		.hps_h2f_lw_axi_master_awid                                        (hps_h2f_lw_axi_master_awid),                              //                                       hps_h2f_lw_axi_master.awid
		.hps_h2f_lw_axi_master_awaddr                                      (hps_h2f_lw_axi_master_awaddr),                            //                                                            .awaddr
		.hps_h2f_lw_axi_master_awlen                                       (hps_h2f_lw_axi_master_awlen),                             //                                                            .awlen
		.hps_h2f_lw_axi_master_awsize                                      (hps_h2f_lw_axi_master_awsize),                            //                                                            .awsize
		.hps_h2f_lw_axi_master_awburst                                     (hps_h2f_lw_axi_master_awburst),                           //                                                            .awburst
		.hps_h2f_lw_axi_master_awlock                                      (hps_h2f_lw_axi_master_awlock),                            //                                                            .awlock
		.hps_h2f_lw_axi_master_awcache                                     (hps_h2f_lw_axi_master_awcache),                           //                                                            .awcache
		.hps_h2f_lw_axi_master_awprot                                      (hps_h2f_lw_axi_master_awprot),                            //                                                            .awprot
		.hps_h2f_lw_axi_master_awvalid                                     (hps_h2f_lw_axi_master_awvalid),                           //                                                            .awvalid
		.hps_h2f_lw_axi_master_awready                                     (hps_h2f_lw_axi_master_awready),                           //                                                            .awready
		.hps_h2f_lw_axi_master_wid                                         (hps_h2f_lw_axi_master_wid),                               //                                                            .wid
		.hps_h2f_lw_axi_master_wdata                                       (hps_h2f_lw_axi_master_wdata),                             //                                                            .wdata
		.hps_h2f_lw_axi_master_wstrb                                       (hps_h2f_lw_axi_master_wstrb),                             //                                                            .wstrb
		.hps_h2f_lw_axi_master_wlast                                       (hps_h2f_lw_axi_master_wlast),                             //                                                            .wlast
		.hps_h2f_lw_axi_master_wvalid                                      (hps_h2f_lw_axi_master_wvalid),                            //                                                            .wvalid
		.hps_h2f_lw_axi_master_wready                                      (hps_h2f_lw_axi_master_wready),                            //                                                            .wready
		.hps_h2f_lw_axi_master_bid                                         (hps_h2f_lw_axi_master_bid),                               //                                                            .bid
		.hps_h2f_lw_axi_master_bresp                                       (hps_h2f_lw_axi_master_bresp),                             //                                                            .bresp
		.hps_h2f_lw_axi_master_bvalid                                      (hps_h2f_lw_axi_master_bvalid),                            //                                                            .bvalid
		.hps_h2f_lw_axi_master_bready                                      (hps_h2f_lw_axi_master_bready),                            //                                                            .bready
		.hps_h2f_lw_axi_master_arid                                        (hps_h2f_lw_axi_master_arid),                              //                                                            .arid
		.hps_h2f_lw_axi_master_araddr                                      (hps_h2f_lw_axi_master_araddr),                            //                                                            .araddr
		.hps_h2f_lw_axi_master_arlen                                       (hps_h2f_lw_axi_master_arlen),                             //                                                            .arlen
		.hps_h2f_lw_axi_master_arsize                                      (hps_h2f_lw_axi_master_arsize),                            //                                                            .arsize
		.hps_h2f_lw_axi_master_arburst                                     (hps_h2f_lw_axi_master_arburst),                           //                                                            .arburst
		.hps_h2f_lw_axi_master_arlock                                      (hps_h2f_lw_axi_master_arlock),                            //                                                            .arlock
		.hps_h2f_lw_axi_master_arcache                                     (hps_h2f_lw_axi_master_arcache),                           //                                                            .arcache
		.hps_h2f_lw_axi_master_arprot                                      (hps_h2f_lw_axi_master_arprot),                            //                                                            .arprot
		.hps_h2f_lw_axi_master_arvalid                                     (hps_h2f_lw_axi_master_arvalid),                           //                                                            .arvalid
		.hps_h2f_lw_axi_master_arready                                     (hps_h2f_lw_axi_master_arready),                           //                                                            .arready
		.hps_h2f_lw_axi_master_rid                                         (hps_h2f_lw_axi_master_rid),                               //                                                            .rid
		.hps_h2f_lw_axi_master_rdata                                       (hps_h2f_lw_axi_master_rdata),                             //                                                            .rdata
		.hps_h2f_lw_axi_master_rresp                                       (hps_h2f_lw_axi_master_rresp),                             //                                                            .rresp
		.hps_h2f_lw_axi_master_rlast                                       (hps_h2f_lw_axi_master_rlast),                             //                                                            .rlast
		.hps_h2f_lw_axi_master_rvalid                                      (hps_h2f_lw_axi_master_rvalid),                            //                                                            .rvalid
		.hps_h2f_lw_axi_master_rready                                      (hps_h2f_lw_axi_master_rready),                            //                                                            .rready
		.config_clk_out_clk_clk                                            (config_clk_clk),                                          //                                          config_clk_out_clk.clk
		.hps_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_003_reset_out_reset),                      // hps_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.pipe_stage_host_ctrl_reset_reset_bridge_in_reset_reset            (rst_controller_reset_out_reset),                          //            pipe_stage_host_ctrl_reset_reset_bridge_in_reset.reset
		.pipe_stage_host_ctrl_s0_address                                   (mm_interconnect_1_pipe_stage_host_ctrl_s0_address),       //                                     pipe_stage_host_ctrl_s0.address
		.pipe_stage_host_ctrl_s0_write                                     (mm_interconnect_1_pipe_stage_host_ctrl_s0_write),         //                                                            .write
		.pipe_stage_host_ctrl_s0_read                                      (mm_interconnect_1_pipe_stage_host_ctrl_s0_read),          //                                                            .read
		.pipe_stage_host_ctrl_s0_readdata                                  (mm_interconnect_1_pipe_stage_host_ctrl_s0_readdata),      //                                                            .readdata
		.pipe_stage_host_ctrl_s0_writedata                                 (mm_interconnect_1_pipe_stage_host_ctrl_s0_writedata),     //                                                            .writedata
		.pipe_stage_host_ctrl_s0_burstcount                                (mm_interconnect_1_pipe_stage_host_ctrl_s0_burstcount),    //                                                            .burstcount
		.pipe_stage_host_ctrl_s0_byteenable                                (mm_interconnect_1_pipe_stage_host_ctrl_s0_byteenable),    //                                                            .byteenable
		.pipe_stage_host_ctrl_s0_readdatavalid                             (mm_interconnect_1_pipe_stage_host_ctrl_s0_readdatavalid), //                                                            .readdatavalid
		.pipe_stage_host_ctrl_s0_waitrequest                               (mm_interconnect_1_pipe_stage_host_ctrl_s0_waitrequest),   //                                                            .waitrequest
		.pipe_stage_host_ctrl_s0_debugaccess                               (mm_interconnect_1_pipe_stage_host_ctrl_s0_debugaccess)    //                                                            .debugaccess
	);

	system_acl_iface_mm_interconnect_2 mm_interconnect_2 (
		.config_clk_out_clk_clk                                 (config_clk_clk),                                            //                               config_clk_out_clk.clk
		.pipe_stage_host_ctrl_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                            // pipe_stage_host_ctrl_reset_reset_bridge_in_reset.reset
		.pipe_stage_host_ctrl_m0_address                        (pipe_stage_host_ctrl_m0_address),                           //                          pipe_stage_host_ctrl_m0.address
		.pipe_stage_host_ctrl_m0_waitrequest                    (pipe_stage_host_ctrl_m0_waitrequest),                       //                                                 .waitrequest
		.pipe_stage_host_ctrl_m0_burstcount                     (pipe_stage_host_ctrl_m0_burstcount),                        //                                                 .burstcount
		.pipe_stage_host_ctrl_m0_byteenable                     (pipe_stage_host_ctrl_m0_byteenable),                        //                                                 .byteenable
		.pipe_stage_host_ctrl_m0_read                           (pipe_stage_host_ctrl_m0_read),                              //                                                 .read
		.pipe_stage_host_ctrl_m0_readdata                       (pipe_stage_host_ctrl_m0_readdata),                          //                                                 .readdata
		.pipe_stage_host_ctrl_m0_readdatavalid                  (pipe_stage_host_ctrl_m0_readdatavalid),                     //                                                 .readdatavalid
		.pipe_stage_host_ctrl_m0_write                          (pipe_stage_host_ctrl_m0_write),                             //                                                 .write
		.pipe_stage_host_ctrl_m0_writedata                      (pipe_stage_host_ctrl_m0_writedata),                         //                                                 .writedata
		.pipe_stage_host_ctrl_m0_debugaccess                    (pipe_stage_host_ctrl_m0_debugaccess),                       //                                                 .debugaccess
		.acl_kernel_interface_ctrl_address                      (mm_interconnect_2_acl_kernel_interface_ctrl_address),       //                        acl_kernel_interface_ctrl.address
		.acl_kernel_interface_ctrl_write                        (mm_interconnect_2_acl_kernel_interface_ctrl_write),         //                                                 .write
		.acl_kernel_interface_ctrl_read                         (mm_interconnect_2_acl_kernel_interface_ctrl_read),          //                                                 .read
		.acl_kernel_interface_ctrl_readdata                     (mm_interconnect_2_acl_kernel_interface_ctrl_readdata),      //                                                 .readdata
		.acl_kernel_interface_ctrl_writedata                    (mm_interconnect_2_acl_kernel_interface_ctrl_writedata),     //                                                 .writedata
		.acl_kernel_interface_ctrl_burstcount                   (mm_interconnect_2_acl_kernel_interface_ctrl_burstcount),    //                                                 .burstcount
		.acl_kernel_interface_ctrl_byteenable                   (mm_interconnect_2_acl_kernel_interface_ctrl_byteenable),    //                                                 .byteenable
		.acl_kernel_interface_ctrl_readdatavalid                (mm_interconnect_2_acl_kernel_interface_ctrl_readdatavalid), //                                                 .readdatavalid
		.acl_kernel_interface_ctrl_waitrequest                  (mm_interconnect_2_acl_kernel_interface_ctrl_waitrequest),   //                                                 .waitrequest
		.acl_kernel_interface_ctrl_debugaccess                  (mm_interconnect_2_acl_kernel_interface_ctrl_debugaccess),   //                                                 .debugaccess
		.version_id_s_read                                      (mm_interconnect_2_version_id_s_read),                       //                                     version_id_s.read
		.version_id_s_readdata                                  (mm_interconnect_2_version_id_s_readdata)                    //                                                 .readdata
	);

	system_acl_iface_mm_interconnect_3 mm_interconnect_3 (
		.pll_outclk0_clk                                              (pll_outclk0_clk),                                                             //                                            pll_outclk0.clk
		.clock_cross_kernel_mem1_m0_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                                          // clock_cross_kernel_mem1_m0_reset_reset_bridge_in_reset.reset
		.clock_cross_kernel_mem1_m0_address                           (clock_cross_kernel_mem1_m0_address),                                          //                             clock_cross_kernel_mem1_m0.address
		.clock_cross_kernel_mem1_m0_waitrequest                       (clock_cross_kernel_mem1_m0_waitrequest),                                      //                                                       .waitrequest
		.clock_cross_kernel_mem1_m0_burstcount                        (clock_cross_kernel_mem1_m0_burstcount),                                       //                                                       .burstcount
		.clock_cross_kernel_mem1_m0_byteenable                        (clock_cross_kernel_mem1_m0_byteenable),                                       //                                                       .byteenable
		.clock_cross_kernel_mem1_m0_read                              (clock_cross_kernel_mem1_m0_read),                                             //                                                       .read
		.clock_cross_kernel_mem1_m0_readdata                          (clock_cross_kernel_mem1_m0_readdata),                                         //                                                       .readdata
		.clock_cross_kernel_mem1_m0_readdatavalid                     (clock_cross_kernel_mem1_m0_readdatavalid),                                    //                                                       .readdatavalid
		.clock_cross_kernel_mem1_m0_write                             (clock_cross_kernel_mem1_m0_write),                                            //                                                       .write
		.clock_cross_kernel_mem1_m0_writedata                         (clock_cross_kernel_mem1_m0_writedata),                                        //                                                       .writedata
		.clock_cross_kernel_mem1_m0_debugaccess                       (clock_cross_kernel_mem1_m0_debugaccess),                                      //                                                       .debugaccess
		.address_span_extender_kernel_windowed_slave_address          (mm_interconnect_3_address_span_extender_kernel_windowed_slave_address),       //            address_span_extender_kernel_windowed_slave.address
		.address_span_extender_kernel_windowed_slave_write            (mm_interconnect_3_address_span_extender_kernel_windowed_slave_write),         //                                                       .write
		.address_span_extender_kernel_windowed_slave_read             (mm_interconnect_3_address_span_extender_kernel_windowed_slave_read),          //                                                       .read
		.address_span_extender_kernel_windowed_slave_readdata         (mm_interconnect_3_address_span_extender_kernel_windowed_slave_readdata),      //                                                       .readdata
		.address_span_extender_kernel_windowed_slave_writedata        (mm_interconnect_3_address_span_extender_kernel_windowed_slave_writedata),     //                                                       .writedata
		.address_span_extender_kernel_windowed_slave_burstcount       (mm_interconnect_3_address_span_extender_kernel_windowed_slave_burstcount),    //                                                       .burstcount
		.address_span_extender_kernel_windowed_slave_byteenable       (mm_interconnect_3_address_span_extender_kernel_windowed_slave_byteenable),    //                                                       .byteenable
		.address_span_extender_kernel_windowed_slave_readdatavalid    (mm_interconnect_3_address_span_extender_kernel_windowed_slave_readdatavalid), //                                                       .readdatavalid
		.address_span_extender_kernel_windowed_slave_waitrequest      (mm_interconnect_3_address_span_extender_kernel_windowed_slave_waitrequest)    //                                                       .waitrequest
	);

	system_acl_iface_irq_mapper irq_mapper (
		.clk           (),                         //       clk.clk
		.reset         (),                         // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq), // receiver0.irq
		.sender_irq    (hps_f2h_irq0_irq)          //    sender.irq
	);

	system_acl_iface_irq_mapper_001 irq_mapper_001 (
		.clk        (),                 //       clk.clk
		.reset      (),                 // clk_reset.reset
		.sender_irq (hps_f2h_irq1_irq)  //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_n),                       // reset_in0.reset
		.clk            (config_clk_clk),                 //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~acl_kernel_interface_sw_reset_export_reset), // reset_in0.reset
		.clk            (pll_outclk0_clk),                             //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),          // reset_out.reset
		.reset_req      (),                                            // (terminated)
		.reset_req_in0  (1'b0),                                        // (terminated)
		.reset_in1      (1'b0),                                        // (terminated)
		.reset_req_in1  (1'b0),                                        // (terminated)
		.reset_in2      (1'b0),                                        // (terminated)
		.reset_req_in2  (1'b0),                                        // (terminated)
		.reset_in3      (1'b0),                                        // (terminated)
		.reset_req_in3  (1'b0),                                        // (terminated)
		.reset_in4      (1'b0),                                        // (terminated)
		.reset_req_in4  (1'b0),                                        // (terminated)
		.reset_in5      (1'b0),                                        // (terminated)
		.reset_req_in5  (1'b0),                                        // (terminated)
		.reset_in6      (1'b0),                                        // (terminated)
		.reset_req_in6  (1'b0),                                        // (terminated)
		.reset_in7      (1'b0),                                        // (terminated)
		.reset_req_in7  (1'b0),                                        // (terminated)
		.reset_in8      (1'b0),                                        // (terminated)
		.reset_req_in8  (1'b0),                                        // (terminated)
		.reset_in9      (1'b0),                                        // (terminated)
		.reset_req_in9  (1'b0),                                        // (terminated)
		.reset_in10     (1'b0),                                        // (terminated)
		.reset_req_in10 (1'b0),                                        // (terminated)
		.reset_in11     (1'b0),                                        // (terminated)
		.reset_req_in11 (1'b0),                                        // (terminated)
		.reset_in12     (1'b0),                                        // (terminated)
		.reset_req_in12 (1'b0),                                        // (terminated)
		.reset_in13     (1'b0),                                        // (terminated)
		.reset_req_in13 (1'b0),                                        // (terminated)
		.reset_in14     (1'b0),                                        // (terminated)
		.reset_req_in14 (1'b0),                                        // (terminated)
		.reset_in15     (1'b0),                                        // (terminated)
		.reset_req_in15 (1'b0)                                         // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~hps_h2f_reset_reset),               // reset_in0.reset
		.clk            (pll_outclk0_clk),                    //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (~hps_h2f_reset_reset),               // reset_in0.reset
		.clk            (config_clk_clk),                     //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	assign kernel_clk_snoop_clk = kernel_clk_clk;

endmodule
